module Decoder_tb;
    
endmodule